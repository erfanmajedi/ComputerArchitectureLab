library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mealy_sequence_detector is
    Port ( A : in  STD_LOGIC;
           Clk : in  STD_LOGIC;
           Reset : in  STD_LOGIC;
           B : out  STD_LOGIC);
end mealy_sequence_detector;

architecture Behavioral of mealy_sequence_detector is
	type state is (s0, s1, s2, s3);
	signal present_state, next_state : state := s0;
	
begin
	syncronous_process : process (clk)
	begin
		if rising_edge(clk) then
			if (Reset = '0') then
				present_state <= s0;
			else
				present_state <= next_state;
			end if;
		end if;
	end process;
 
	next_state_and_output_decoder : process(present_state, A)
	begin
		B <= '0'; 
		case (present_state) is 
			when s0 =>
				if (A = '1') then
					next_state <= s1;
					B <= '0';
				else
					next_state <= s0;
					B <= '0'; 
				end if; 
			when s1 =>
				if (A = '1') then
					next_state <= s2;
					B <= '0';
				else
					next_state <= s0;
					B <= '0'; 
				end if; 
			when s2 =>
				if (A = '1') then
					next_state <= s2;
					B <= '0';
				else
					next_state <= s3;
					B <= '0'; 
				end if; 
			when s3 =>
				if (A = '1') then
					next_state <= s2;
					B <= '1';
				else
					next_state <= s0;
					B <= '0'; 
				end if; 
			when others =>
				next_state <= s0;
				B <= '0';
		end case;
	end process;
end Behavioral;

